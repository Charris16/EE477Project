../../verilog/opcode.vh